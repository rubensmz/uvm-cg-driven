class cg_driven_subscriber extends uvm_subscriber;

endclass : cg_driven_subscriber