module dut(input [3:0] addr, data, input clk);

endmodule