class cg_subscriber extends uvm_subscriber;

endclass : cg_subscriber