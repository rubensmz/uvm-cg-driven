interface pkt_if;
    logic [3:0] addr;
    logic [3:0] data;
endinterface : pkt_if