package cg_driven_pkg;
    `include "uvm_macros.svh"
    import uvm_pkg::*;

    import pkt_agent_pkg::*;

    //`include "cg_driven_subscriber.sv"
    `include "cg_driven_env.sv"
    `include "cg_driven_test.sv"

endpackage : cg_driven_pkg