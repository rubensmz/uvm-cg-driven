`include "pkt_if.sv"

package pkt_agt_pkg;
    `include "pkt_tr.sv"
    `include "pkt_driver.sv"
    `include "pkt_sequencer.sv"
    `include "pkt_monitor.sv"
    `include "pkt_agent.sv"
endpackage : pkt_agt_pkg