interface pkt_if;
    logic [3:0] addr;
    logic [7:0] data;
endinterface : pkt_if