interface pkt_if;
    logic [3:0] addr;
    logic [3:0] data;
    logic clk;
endinterface : pkt_if